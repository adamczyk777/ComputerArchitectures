--karta graficzna w VHDL
